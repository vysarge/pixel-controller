`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/05/2016 09:17:09 AM
// Design Name: 
// Module Name: pattern_modifier
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module pattern_modifier(
    input init,
    input fclock,
    input cclock,
    input [3:0] xin,
    input [3:0] yin,
    input [4:0] rgbin,
    input [3:0] xout,
    input [3:0] yout,
    input [4:0] rgbout
    );
endmodule
